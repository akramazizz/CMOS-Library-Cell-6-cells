*** SPICE deck for cell size1_sim{sch} from library complex_function_1
*** Created on Sun May 16, 2021 18:06:33
*** Last revised on Sun May 16, 2021 18:25:28
*** Written on Mon May 17, 2021 00:54:10 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT complex_function_1__size1 FROM CELL complex_function_1:size1{sch}
.SUBCKT complex_function_1__size1 out w x y z
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@14 y gnd gnd N L=0.2U W=0.8U
Mnmos@1 out x net@14 gnd N L=0.2U W=0.8U
Mnmos@2 out w net@48 gnd N L=0.2U W=0.8U
Mnmos@4 net@48 z gnd gnd N L=0.2U W=0.8U
Mpmos@0 net@8 w out vdd P L=0.2U W=1.952U
Mpmos@1 vdd y net@8 vdd P L=0.2U W=1.952U
Mpmos@2 net@8 z out vdd P L=0.2U W=1.952U
Mpmos@3 vdd x net@8 vdd P L=0.2U W=1.952U
.ENDS complex_function_1__size1

.global gnd vdd

*** TOP LEVEL CELL: complex_function_1:size1_sim{sch}
Xsize1@0 y vdd gnd gnd in complex_function_1__size1

* Spice Code nodes in cell cell 'complex_function_1:size1_sim{sch}'
vdd vdd 0 dc 1.8
vin in 0 DC pulse 0 1.8 0.1n 0p 0p 5n 10n
.tran 0 200n
cload y 0 100fF
.measure tpdr_0_cinv v(in) val=0.9 fall=1 TARG v(y) val=0.9 rise=1
.measure tpdf_0_cinv v(in) val=0.9 rise=1 TARG v(y) val=0.9 fall=1
.include c:\electric\scmos.txt
.END
